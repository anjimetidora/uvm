//***************************************************************************//
//***************************************************************************//
//***************************************************************************//
//**************                                          *******************//
//**************                                          *******************//
//**************      (c) SASIC Technologies Pvt Ltd      *******************//
//**************          (c) Verilogic Solutions         *******************//
//**************                                          *******************//
//**************                                          *******************//
//**************                                          *******************//
//**************           www.sasictek.com               *******************//
//**************          www.verilog-ic.com              *******************//
//**************                                          *******************//
//**************           Twitter:@sasictek              *******************//
//**************                                          *******************//
//**************                                          *******************//
//**************                                          *******************//
//***************************************************************************//
//***************************************************************************//


//              File Name : fifo_sequencer.sv
//              File Type: System Verilog                                 
//              Creation Date : 09-08-2017
//              Last Modified : Wed 09 Aug 2017 10:39:59 AM IST

                             
//***************************************************************************//
//***************************************************************************//
                             

//              Author:
//              Reviewer:
//              Manager:
                             

//***************************************************************************//
//***************************************************************************//


class fifo_sequencer extends uvm_sequencer#(fifo_sequence_item)
`uvm_component_utils(fifo_sequencer)

function new(string name="fifo_sequencer",uvm_component parent)
	begin
		super.new(name,parent);
	end
endfunction

endclass


