//***************************************************************************//
//***************************************************************************//
//***************************************************************************//
//**************                                          *******************//
//**************                                          *******************//
//**************      (c) SASIC Technologies Pvt Ltd      *******************//
//**************          (c) Verilogic Solutions         *******************//
//**************                                          *******************//
//**************                                          *******************//
//**************                                          *******************//
//**************           www.sasictek.com               *******************//
//**************          www.verilog-ic.com              *******************//
//**************                                          *******************//
//**************           Twitter:@sasictek              *******************//
//**************                                          *******************//
//**************                                          *******************//
//**************                                          *******************//
//***************************************************************************//
//***************************************************************************//


//              File Name : fifo_top.sv
//              File Type: System Verilog                                 
//              Creation Date : 09-08-2017
//              Last Modified : Fri 11 Aug 2017 03:30:27 PM IST

                             
//***************************************************************************//
//***************************************************************************//
                             

//              Author:
//              Reviewer:
//              Manager:
                             

//***************************************************************************//
//***************************************************************************//



module fifo_top;

fifo_interface top_inf(.in_clk(top_clk));
	
fifo dut_insta(.rst_n(top_inf.rst_n),
								.push(top_inf.push),
								.pop(top_inf.pop),
								.in_data(top_inf.in_data),
								.data_out(top_inf.data_out),
								.full(top_inf.full),
								.empty(top_inf.empty),
								.push_err_on_full(top_inf.push_err_on_full),
								.pop_err_on_empty(top_inf.pop_err_on_empty));

	
	initial 
		begin
			top_clk='b0;
			forever #5 top_clk=~top_clk;
		end
	
	initial
		begin
			uvm_config_db#(virtual fifo_interface)::set(.cntxt(null),
																									.inst_name("*"),
																									.field_name("top_inf"),
																									.value(top_inf));
			run_test();
		end

endmodule
