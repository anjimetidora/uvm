library verilog;
use verilog.vl_types.all;
entity mc_package is
end mc_package;
