//***************************************************************************//
//***************************************************************************//
//***************************************************************************//
//**************                                          *******************//
//**************                                          *******************//
//**************      (c) SASIC Technologies Pvt Ltd      *******************//
//**************          (c) Verilogic Solutions         *******************//
//**************                                          *******************//
//**************                                          *******************//
//**************                                          *******************//
//**************           www.sasictek.com               *******************//
//**************          www.verilog-ic.com              *******************//
//**************                                          *******************//
//**************           Twitter:@sasictek              *******************//
//**************                                          *******************//
//**************                                          *******************//
//**************                                          *******************//
//***************************************************************************//
//***************************************************************************//


//              File Name : ahbl_package.sv
//              File Type: System Verilog                                 
//              Creation Date : 18-12-2017
//              Last Modified : Mon 18 Dec 2017 12:06:02 PM IST

                             
//***************************************************************************//
//***************************************************************************//
                             

//              Author:
//              Reviewer:
//              Manager:
                             

//***************************************************************************//
//***************************************************************************//


package ahbl_package;

parameter ADDR_WIDTH=32;
parameter SIZE_WIDTH=3;
parameter BURST_WIDTH=3;
parameter PROT_WIDTH=4;
parameter TRANS_WIDTH=2;
parameter WDATA_WIDTH=32;
parameter RDATA_WIDTH=32;

endpackage
