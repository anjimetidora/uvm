//***************************************************************************//
//***************************************************************************//
//***************************************************************************//
//**************                                          *******************//
//**************                                          *******************//
//**************      (c) SASIC Technologies Pvt Ltd      *******************//
//**************          (c) Verilogic Solutions         *******************//
//**************                                          *******************//
//**************                                          *******************//
//**************                                          *******************//
//**************           www.sasictek.com               *******************//
//**************          www.verilog-ic.com              *******************//
//**************                                          *******************//
//**************           Twitter:@sasictek              *******************//
//**************                                          *******************//
//**************                                          *******************//
//**************                                          *******************//
//***************************************************************************//
//***************************************************************************//


//              File Name : ahbl_sequence.sv
//              File Type: System Verilog                                 
//              Creation Date : 18-12-2017
//              Last Modified : Mon 18 Dec 2017 01:02:00 PM IST

                             
//***************************************************************************//
//***************************************************************************//
                             

//              Author:
//              Reviewer:
//              Manager:
                             

//***************************************************************************//
//***************************************************************************//


class ahbl_sequence extends uvm_sequence #(ahbl_sequence_item);
//factory registration
`uvm_object_utils(ahbl_sequence)

function new(string name="ahbl_sequence");
super.new(name);
endfunction

extern virtual task body();

endclass:ahbl_sequence


task ahbl_sequence::body();
`uvm_info(get_name(),$sformatf("sequence is running...........\n"),UVM_LOW)


`uvm_do(req)



`uvm_info(get_name(),$sformatf("sequence is end..............\n"),UVM_LOW)

endtask:task_body




