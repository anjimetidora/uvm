//***************************************************************************//
//***************************************************************************//
//***************************************************************************//
//**************                                          *******************//
//**************                                          *******************//
//**************      (c) SASIC Technologies Pvt Ltd      *******************//
//**************          (c) Verilogic Solutions         *******************//
//**************                                          *******************//
//**************                                          *******************//
//**************                                          *******************//
//**************           www.sasictek.com               *******************//
//**************          www.verilog-ic.com              *******************//
//**************                                          *******************//
//**************           Twitter:@sasictek              *******************//
//**************                                          *******************//
//**************                                          *******************//
//**************                                          *******************//
//***************************************************************************//
//***************************************************************************//


//              File Name : ahbl_sequencer.sv
//              File Type: System Verilog                                 
//              Creation Date : 20-12-2017
//              Last Modified : Wed 20 Dec 2017 01:18:44 PM IST

                             
//***************************************************************************//
//***************************************************************************//
                             

//              Author:
//              Reviewer:
//              Manager:
                             

//***************************************************************************//
//***************************************************************************//

class ahbl_sequencer extends uvm_sequencer #(ahbl_sequence_item)

	`uvm_component_utils(ahbl_sequencer)

	function new(string name="ahbl_sequencer", uvm_component parent);
	super.new(name,parent);
	endfunction
endclass
