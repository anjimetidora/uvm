
`include "read_test/mc_read_seq.sv"
`include "write_test/mc_write_seq.sv"
