//*******************************DV_logic*************************************//

//												File Name : slv_err_seq.sv
//												File Type : system_verilog
//										Creation Date : 26-10-2018
//												File Type : system_verilog
//													 Author : Dorababu

//****************************************************************************//
