//***************************************************************************//
//***************************************************************************//
//***************************************************************************//
//**************                                          *******************//
//**************                                          *******************//
//**************      (c) SASIC Technologies Pvt Ltd      *******************//
//**************          (c) Verilogic Solutions         *******************//
//**************                                          *******************//
//**************                                          *******************//
//**************                                          *******************//
//**************           www.sasictek.com               *******************//
//**************          www.verilog-ic.com              *******************//
//**************                                          *******************//
//**************           Twitter:@sasictek              *******************//
//**************                                          *******************//
//**************                                          *******************//
//**************                                          *******************//
//***************************************************************************//
//***************************************************************************//


//              File Name : ahbl_interface.sv
//              File Type: System Verilog                                 
//              Creation Date : 18-12-2017
//              Last Modified : Mon 18 Dec 2017 12:31:58 PM IST

                             
//***************************************************************************//
//***************************************************************************//
                             

//              Author:
//              Reviewer:
//              Manager:
                             

//***************************************************************************//
//***************************************************************************//
import ahbl_package::*;

interface ahbl_interface #(HCLK);

logic HRESETn;
logic HCLK;
logic [ADDR_WIDTH-1:0]HADDR;
logic HWRITE;
logic [WDATA_WIDTH-1:0]HWDATA;
logic [SIZE_WIDTH-1:0]HSIZE;
logic [BURST_WIDTH-1:0]HBURST;
logic [TRANS_WIDTH-1:0]HTRANS;
logic [PROT_WIDTH-1:0]HPROT;
logic HMAST_LOCK;
logic  HREADY;
logic  HRESP;

clocking drv_cb@(negedge HCLK);
endclocking 

clocking mon_cb@(negedge HCLK);
endclocking

endinterface



