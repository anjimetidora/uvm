package mc_package;

  parameter DATA_WIDTH='d8;
  parameter ADDR_WIDTH='d256;
endpackage


